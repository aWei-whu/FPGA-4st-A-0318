
`timescale 1 ns / 1 ps

  module DownSample_mul_mucud_DSP48_0(a, b, p);
input [6 - 1 : 0] a;
input signed [10 - 1 : 0] b;
output signed [10 - 1 : 0] p;

assign p = $signed ({1'b0, a}) * $signed (b);

endmodule
`timescale 1 ns / 1 ps
module DownSample_mul_mucud(
    din0,
    din1,
    dout);

parameter ID = 32'd1;
parameter NUM_STAGE = 32'd1;
parameter din0_WIDTH = 32'd1;
parameter din1_WIDTH = 32'd1;
parameter dout_WIDTH = 32'd1;
input[din0_WIDTH - 1:0] din0;
input[din1_WIDTH - 1:0] din1;
output[dout_WIDTH - 1:0] dout;



DownSample_mul_mucud_DSP48_0 DownSample_mul_mucud_DSP48_0_U(
    .a( din0 ),
    .b( din1 ),
    .p( dout ));

endmodule

